---------------------------------------------------------------------
-- DEV		: 
-- ACADEMIC : KULEUVEN 2019-2020 CAMPUS DE NAYER
-- MODULE	: 
-- INFO		:  
---------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity "MODULE NAME HERE" is
    port( 
            
    );
end "MODULE NAME HERE";

architecture Behavioral OF "MODULE NAME HERE" IS
-- SIGNALS HERE
begin
-- SYNC COMPONENT HERE

-- COMB COMPONENT HERE

-- LINKING SIGNALS HERE

end Behavioral;
